library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity memory is
  PORT (
    --clka : IN STD_LOGIC;
    wea : IN STD_LOGIC;
    clk : IN std_logic;
    addra : IN STD_LOGIC_VECTOR(0 to 7);
    dina : IN STD_LOGIC_VECTOR(0 to 7);
   -- clkb : IN STD_LOGIC;
    reset : IN std_logic;
    enb : IN STD_LOGIC;
    addrb : IN STD_LOGIC_VECTOR(0 to 7);
    doutb : OUT STD_LOGIC_VECTOR(0 to 7)
  );
end memory;

architecture Behavioral of memory is

	type Memory_type is array (0 to 255) of std_logic_vector (0 to 7);
	signal Memory_array : Memory_type;
	signal manoj : Memory_type;
	signal address : unsigned (0 to 7);
	signal clka : std_logic;
	signal clkb : std_logic;
	signal temp : integer;
	signal temp1 : integer;
	
begin

process(clk)
    begin
        if(clk'event and clk = '1') then
        temp <= temp+1;
        if(temp = 325) then
            clka <= not clka;
            temp <= 0;
        end if;
      end if;
end process;

    process(clk, reset)
    begin
    if(reset = '1') then
        temp1 <= 0;
            elsif(clk'event and clk = '1') then
        temp1 <= temp1+1;
        if(temp1 = 5208) then
            clkb <= not clkb;
            temp1 <= 0;
        end if;
      end if;
    end process;

--    process( clkb)
--    begin
--      if(reset = '1') then
--        doutb <= "00000000";
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  
--      end if;
--    end process;

	process (clkb)
	begin
    if rising_edge(clkb) then    
        if (enb = '1') then
            address <= unsigned(addrb);    
        end if;
    end if;
    end process;
	doutb <= Memory_array (to_integer(address));
	process (clkb)
	begin
		if rising_edge(clkb) then	
			if (wea = '1') then
				Memory_array (to_integer(unsigned(addra))) <= dina (0 to 7);	
			end if;
		end if;
	end process;
end Behavioral;
